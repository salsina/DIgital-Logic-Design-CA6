module tb();
  reg[15:0] x;
  reg[7:0] y;
  reg start,clk,rst;
  wire ready;
  wire [15:0] sinx;
  datapath dp(x,y,start,clk,rst,sinx, ready);
  initial begin
    rst = 1;
    clk = 0;
    start = 0;
    x = 0000000110001000 ;
    y = 00000001;
    #30 rst = 0;
    start = 1;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
     start = 0;    
    
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;       
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;       
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;       
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;       
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;       
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;           
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;       
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;
    #30 clk = 1;
    #30 clk = 0;       
  end
endmodule